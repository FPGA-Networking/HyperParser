`timescale  1ns / 1ps

module tb_test_pex_ibf_pdep_bf_top;

// test_pex_ibf_pdep_bf_top Parameters
parameter PERIOD      = 10;
parameter DATA_WIDTH  = 4096;



parameter MODE_WIDTH                  = 2; // 2 ,
parameter IBF_CFG_WIDTH_2_2           = DATA_WIDTH/2 ; //单级stage的config width
parameter IBF_N_NUM_2_1               = 32;//32 ,
parameter IBF_CFG_WIDTH_2_1           = $clog2(IBF_N_NUM_2_1)*(DATA_WIDTH/IBF_N_NUM_2_1) ;

parameter BF_CFG_WIDTH_2_2            = (DATA_WIDTH/(2*8))/4 ; // 除4是因为4个segment
                








// test_pex_ibf_pdep_bf_top Inputs
reg   clk                                  = 0 ;
reg   rst                                  = 1 ;
reg   [MODE_WIDTH-1:0]  mode_i             = 0 ;
reg   dval_i                               = 0 ;
reg   [DATA_WIDTH-1:0]  data_i             = 0 ;
reg   [7:0]  ibf_sram_sel_2_2              = 0 ;
reg   ibf_wr_en_2_2                        = 0 ;
reg   [IBF_CFG_WIDTH_2_2-1:0]  ibf_wr_cfg_2_2 = 0 ;
reg   ibf_wr_en_2_1                        = 0 ;
reg   [IBF_CFG_WIDTH_2_1-1:0]  ibf_wr_cfg_2_1 = 0 ;
reg   [7:0]  bf_sram_sel_2_2               = 0 ;
reg   bf_wr_en_2_2_A                         = 0 ;
reg   bf_wr_en_2_2_B                         = 0 ;
reg   bf_wr_en_2_2_C                         = 0 ;
reg   bf_wr_en_2_2_D                         = 0 ;
reg   [BF_CFG_WIDTH_2_2-1:0]  bf_wr_cfg_2_2 = 0 ;

// test_pex_ibf_pdep_bf_top Outputs
wire  dval_o                               ;
wire  [DATA_WIDTH-1:0]  data_o             ;


initial
begin
    forever #(PERIOD/2)  clk=~clk;
end

initial
begin
    #(PERIOD*2) rst  =  0;
end


reg   [MODE_WIDTH-1:0]  mode_temp_1             = 0 ;
reg                     dval_temp_1             = 0 ;
reg   [DATA_WIDTH-1:0]  data_temp_1             = 0 ;

reg   [MODE_WIDTH-1:0]  mode_temp_2             = 0 ;
reg                     dval_temp_2             = 0 ;
reg   [DATA_WIDTH-1:0]  data_temp_2             = 0 ;

reg   [MODE_WIDTH-1:0]  mode_temp_3             = 0 ;
reg                     dval_temp_3             = 0 ;
reg   [DATA_WIDTH-1:0]  data_temp_3             = 0 ;

reg   [MODE_WIDTH-1:0]  mode_temp_4             = 0 ;
reg                     dval_temp_4             = 0 ;
reg   [DATA_WIDTH-1:0]  data_temp_4             = 0 ;

reg   [MODE_WIDTH-1:0]  mode_temp_5             = 0 ;
reg                     dval_temp_5             = 0 ;
reg   [DATA_WIDTH-1:0]  data_temp_5             = 0 ;

reg   [MODE_WIDTH-1:0]  mode_temp_6             = 0 ;
reg                     dval_temp_6             = 0 ;
reg   [DATA_WIDTH-1:0]  data_temp_6             = 0 ;


always @(posedge clk) begin
    mode_temp_1 <=  mode_i ;
    dval_temp_1 <=  dval_i ;
    data_temp_1 <=  data_i ;
    mode_temp_2 <= mode_temp_1 ; 
    dval_temp_2 <= dval_temp_1 ; 
    data_temp_2 <= data_temp_1 ; 
    mode_temp_3 <= mode_temp_2 ; 
    dval_temp_3 <= dval_temp_2 ; 
    data_temp_3 <= data_temp_2 ; 
    mode_temp_4 <= mode_temp_3 ; 
    dval_temp_4 <= dval_temp_3 ; 
    data_temp_4 <= data_temp_3 ; 
    mode_temp_5 <= mode_temp_4 ; 
    dval_temp_5 <= dval_temp_4 ; 
    data_temp_5 <= data_temp_4 ; 
    mode_temp_6 <= mode_temp_5 ; 
    dval_temp_6 <= dval_temp_5 ; 
    data_temp_6 <= data_temp_5 ; 
end



test_pex_ibf_pdep_bf_top u_test_pex_ibf_pdep_bf_top(
    .clk              (clk              ),
    // .rst              (1'b0              ),
    .mode_i           (mode_temp_1           ),
    .dval_i           (dval_temp_3           ),
    .data_i           (data_temp_3           ),
    .dval_o           (dval_o           ),
    .data_o           (data_o           ),
    // .ibf_sram_sel_2_2 (ibf_sram_sel_2_2 ),
    // .ibf_wr_en_2_2    (ibf_wr_en_2_2    ),
    // .ibf_wr_cfg_2_2   (ibf_wr_cfg_2_2   ),
    // .ibf_wr_en_2_1    (ibf_wr_en_2_1    ),
    // .ibf_wr_cfg_2_1   (ibf_wr_cfg_2_1   ),
    // .bf_sram_sel_2_2  (bf_sram_sel_2_2  ),
    // .bf_wr_en_2_2_A     (bf_wr_en_2_2_A     ),
    // .bf_wr_en_2_2_B     (bf_wr_en_2_2_B     ),
    // .bf_wr_en_2_2_C     (bf_wr_en_2_2_C     ),
    // .bf_wr_en_2_2_D     (bf_wr_en_2_2_D     ),

    // .bf_wr_cfg_2_2    (bf_wr_cfg_2_2    ),

    .cfg_sel_module   ( 2'b0 )    ,
    .cfg_sram_sel     ( 8'b0 )    ,
    .cfg_addr_write   ( 7'b0 )    ,
    .cfg_wr_en        ( 1'b0 )    ,
    .cfg_data         ( 64'b0 )        



);






// b1000_0001_0010_1011

// 对于pex，mode=0对应的是提取第二个4bit，mode=1对应的是提取前4个bit的第一个bit，mode=2对应的是提取最后4bit


// 对于pdep，测试了4种模式，[1,1,0,0]，初始值是['3', '0']，[1,0,1,0]与['2', '1']，[0,1,0,1]与['2', '2']，[0,1,1,0]与['2', '3']

initial
begin
// seg 4096    
    #200
    dval_i = 1'b1;
    mode_i  = 2'b00;
    data_i = 4096'heed6640c13fe75b83ed539a90800057ce2d64b9b0000d80105f530670ec2cc88562808d026088e40d32673a2e35fb5b299daed825e965c312173fac60000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//ICMP 提取000100000000010000
    #(PERIOD)
    dval_i = 'b0;
    mode_i  = 2'b00;
    data_i = 'b0;
    #200
    dval_i = 1'b1;
    mode_i  = 2'b00;
    data_i = 4096'h4a73219fbcbeb2f0bc4c0169080006ae718916430000a0062556575a2878d7e1974021e21a3668134f6072ba6624aa7064bd5076a8eabfd309c933a80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//TCP 提取000000000110101000
    #(PERIOD)
    dval_i = 'b0;
    mode_i  = 2'b00;
    data_i = 'b0;
    #200
    dval_i = 1'b1;
    mode_i  = 2'b00;
    data_i = 4096'h5860481e6a3e240908b57e84080005bc2637025b00006c11078364a10cced39c4e31d981000069aa4a541b1f9c153d402051f37b0127e98f20776c8e0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//UDP 提取000010001000000011
    #(PERIOD)
    dval_i = 'b0;
    mode_i  = 2'b00;
    data_i = 'b0;


// seg 2048
    #200
    dval_i = 1'b1;
    mode_i  = 2'b01;
    data_i = 4096'heed6640c13fe75b83ed539a90800057ce2d64b9b0000d80105f530670ec2cc88562808d026088e40d32673a2e35fb5b299daed825e965c312173fac600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000eed6640c13fe75b83ed539a90800057ce2d64b9b0000d80105f530670ec2cc88562808d026088e40d32673a2e35fb5b299daed825e965c312173fac600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//ICMP 提取000100000000010000
    #(PERIOD)
    dval_i = 'b0;
    mode_i  = 2'b00;
    data_i = 'b0;
    #200
    dval_i = 1'b1;
    mode_i  = 2'b01;
    data_i = 4096'h4a73219fbcbeb2f0bc4c0169080006ae718916430000a0062556575a2878d7e1974021e21a3668134f6072ba6624aa7064bd5076a8eabfd309c933a8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004a73219fbcbeb2f0bc4c0169080006ae718916430000a0062556575a2878d7e1974021e21a3668134f6072ba6624aa7064bd5076a8eabfd309c933a800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//TCP 提取000000000110101000
    #(PERIOD)
    dval_i = 'b0;
    mode_i  = 2'b00;
    data_i = 'b0;
    #200
    dval_i = 1'b1;
    mode_i  = 2'b01;
    data_i = 4096'h5860481e6a3e240908b57e84080005bc2637025b00006c11078364a10cced39c4e31d981000069aa4a541b1f9c153d402051f37b0127e98f20776c8e000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005860481e6a3e240908b57e84080005bc2637025b00006c11078364a10cced39c4e31d981000069aa4a541b1f9c153d402051f37b0127e98f20776c8e00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//UDP 提取000010001000000011
    #(PERIOD)
    dval_i = 'b0;
    mode_i  = 2'b00;
    data_i = 'b0;


// seg 1024
    #200
    dval_i = 1'b1;
    mode_i  = 2'b10;
    data_i = 4096'heed6640c13fe75b83ed539a90800057ce2d64b9b0000d80105f530670ec2cc88562808d026088e40d32673a2e35fb5b299daed825e965c312173fac60000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000eed6640c13fe75b83ed539a90800057ce2d64b9b0000d80105f530670ec2cc88562808d026088e40d32673a2e35fb5b299daed825e965c312173fac60000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000eed6640c13fe75b83ed539a90800057ce2d64b9b0000d80105f530670ec2cc88562808d026088e40d32673a2e35fb5b299daed825e965c312173fac60000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000eed6640c13fe75b83ed539a90800057ce2d64b9b0000d80105f530670ec2cc88562808d026088e40d32673a2e35fb5b299daed825e965c312173fac60000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//ICMP 提取000100000000010000
    #(PERIOD)
    dval_i = 'b0;
    mode_i  = 2'b00;
    data_i = 'b0;
    #200
    dval_i = 1'b1;
    mode_i  = 2'b10;
    data_i = 4096'h4a73219fbcbeb2f0bc4c0169080006ae718916430000a0062556575a2878d7e1974021e21a3668134f6072ba6624aa7064bd5076a8eabfd309c933a800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004a73219fbcbeb2f0bc4c0169080006ae718916430000a0062556575a2878d7e1974021e21a3668134f6072ba6624aa7064bd5076a8eabfd309c933a800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004a73219fbcbeb2f0bc4c0169080006ae718916430000a0062556575a2878d7e1974021e21a3668134f6072ba6624aa7064bd5076a8eabfd309c933a800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004a73219fbcbeb2f0bc4c0169080006ae718916430000a0062556575a2878d7e1974021e21a3668134f6072ba6624aa7064bd5076a8eabfd309c933a80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//TCP 提取000000000110101000
    #(PERIOD)
    dval_i = 'b0;
    mode_i  = 2'b00;
    data_i = 'b0;
    #200
    dval_i = 1'b1;
    mode_i  = 2'b10;
    data_i = 4096'h5860481e6a3e240908b57e84080005bc2637025b00006c11078364a10cced39c4e31d981000069aa4a541b1f9c153d402051f37b0127e98f20776c8e00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005860481e6a3e240908b57e84080005bc2637025b00006c11078364a10cced39c4e31d981000069aa4a541b1f9c153d402051f37b0127e98f20776c8e00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005860481e6a3e240908b57e84080005bc2637025b00006c11078364a10cced39c4e31d981000069aa4a541b1f9c153d402051f37b0127e98f20776c8e00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005860481e6a3e240908b57e84080005bc2637025b00006c11078364a10cced39c4e31d981000069aa4a541b1f9c153d402051f37b0127e98f20776c8e0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//UDP 提取000010001000000011
    #(PERIOD)
    dval_i = 'b0;
    mode_i  = 2'b00;
    data_i = 'b0;






















    // #200
    // dval_i = 1'b1;
    // data_i = 16'b1001_0001_0001_1111;
    // #(PERIOD)
    // dval_i = 'b0;
    // data_i = 'b0;
end



// initial
// begin
//     #200
//     dval_i = 1'b1;
//     mode_i  = 2'b00;
//     data_i = 4096'h4a73219fbcbeb2f0bc4c0169080006ae718916430000a0062556575a2878d7e1974021e21a3668134f6072ba6624aa7064bd5076a8eabfd309c933a80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//ICMP 提取000100000000010000
//     #(PERIOD)
//     dval_i = 'b0;
//     mode_i  = 2'b00;
//     data_i = 'b0;
//     #200
//     dval_i = 1'b1;
//     mode_i  = 2'b01;
//     data_i = 4096'h4a73219fbcbeb2f0bc4c0169080006ae718916430000a0062556575a2878d7e1974021e21a3668134f6072ba6624aa7064bd5076a8eabfd309c933a80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//TCP 提取000000000110101000
//     #(PERIOD)
//     dval_i = 'b0;
//     mode_i  = 2'b00;
//     data_i = 'b0;
//     #200
//     dval_i = 1'b1;
//     mode_i  = 2'b10;
//     data_i = 4096'h4a73219fbcbeb2f0bc4c0169080006ae718916430000a0062556575a2878d7e1974021e21a3668134f6072ba6624aa7064bd5076a8eabfd309c933a80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//UDP 提取000010001000000011
//     #(PERIOD)
//     dval_i = 'b0;
//     mode_i  = 2'b00;
//     data_i = 'b0;
//     // #200
//     // dval_i = 1'b1;
//     // data_i = 16'b1001_0001_0001_1111;
//     // #(PERIOD)
//     // dval_i = 'b0;
//     // data_i = 'b0;
// end




parameter ICMP_BIT_MASK_SEG_01 = 4096'hffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
parameter TCP_BIT_MASK_SEG_01  = 4096'hffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
parameter UDP_BIT_MASK_SEG_01  = 4096'hffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffff000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


parameter ICMP_BIT_PHV_SEG_01 = 4096'heed6640c13fe75b83ed539a908000000000000000000057ce2d64b9b0000d80105f530670ec2cc885628000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008d026080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
parameter TCP_BIT_PHV_SEG_01  = 4096'h4a73219fbcbeb2f0bc4c01690800000000000000000006ae718916430000a0062556575a2878d7e197400000000000000000000000000000000000000000000000000000000000000000000000000000000021e21a3668134f6072ba6624aa7064bd5076a8ea0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
parameter UDP_BIT_PHV_SEG_01  = 4096'h5860481e6a3e240908b57e840800000000000000000005bc2637025b00006c11078364a10cced39c4e31000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d981000069aa4a54000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


reg result_correct_SEG_01 = 1'b0 ;
reg [4095:0] data_temp_icmp_SEG_01 = 'b0 ;
reg [4095:0] data_temp_tcp_SEG_01  = 'b0 ;
reg [4095:0] data_temp_udp_SEG_01  = 'b0 ;
wire [4095:0] wire_data_temp_icmp_SEG_01  ;
wire [4095:0] wire_data_temp_tcp_SEG_01   ;
wire [4095:0] wire_data_temp_udp_SEG_01   ;


assign wire_data_temp_icmp_SEG_01 =  data_o&ICMP_BIT_MASK_SEG_01;
assign wire_data_temp_tcp_SEG_01  =  data_o&TCP_BIT_MASK_SEG_01;
assign wire_data_temp_udp_SEG_01  =  data_o&UDP_BIT_MASK_SEG_01;

reg flag_icmp_SEG_01 ;
reg flag_tcp_SEG_01  ;
reg flag_udp_SEG_01  ;

always @(negedge clk) begin
    // if ( dval_o == 1'b1 ) begin
        data_temp_icmp_SEG_01 <= (data_o&ICMP_BIT_MASK_SEG_01)^ICMP_BIT_PHV_SEG_01    ;
        data_temp_tcp_SEG_01  <= (data_o&TCP_BIT_MASK_SEG_01 )^TCP_BIT_PHV_SEG_01     ;
        data_temp_udp_SEG_01  <= (data_o&UDP_BIT_MASK_SEG_01 )^UDP_BIT_PHV_SEG_01     ;
        
        flag_icmp_SEG_01 <=  ((data_o&ICMP_BIT_MASK_SEG_01) == ICMP_BIT_PHV_SEG_01); // |((data_o&ICMP_BIT_MASK)^ICMP_BIT_PHV ) ;
        flag_tcp_SEG_01  <= |((data_o&TCP_BIT_MASK_SEG_01 )^TCP_BIT_PHV_SEG_01  ) ;
        flag_udp_SEG_01  <= |((data_o&UDP_BIT_MASK_SEG_01 )^UDP_BIT_PHV_SEG_01  ) ;


        if ( !((data_o&ICMP_BIT_MASK_SEG_01)^ICMP_BIT_PHV_SEG_01) ) begin // data_o&ICMP_BIT_MASK == ICMP_BIT_PHV
            result_correct_SEG_01 <= 1'b1;
        end
        else if (!((data_o&TCP_BIT_MASK_SEG_01 )^TCP_BIT_PHV_SEG_01)) begin // data_o&TCP_BIT_MASK == TCP_BIT_PHV
            result_correct_SEG_01 <= 1'b1;
        end
        else if(!((data_o&UDP_BIT_MASK_SEG_01 )^UDP_BIT_PHV_SEG_01)) begin // data_o&UDP_BIT_MASK == UDP_BIT_PHV
            result_correct_SEG_01 <= 1'b1;
        end
        else begin
            result_correct_SEG_01 <= 1'b0;
        end
    // end
end




parameter ICMP_BIT_MASK_SEG_02 = 4096'hffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
parameter TCP_BIT_MASK_SEG_02  = 4096'hffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
parameter UDP_BIT_MASK_SEG_02  = 4096'hffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


parameter ICMP_BIT_PHV_SEG_02 = 4096'heed6640c13fe75b83ed539a908000000000000000000057ce2d64b9b0000d80105f530670ec2cc885628000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008d0260800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000eed6640c13fe75b83ed539a908000000000000000000057ce2d64b9b0000d80105f530670ec2cc885628000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008d0260800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
parameter TCP_BIT_PHV_SEG_02  = 4096'h4a73219fbcbeb2f0bc4c01690800000000000000000006ae718916430000a0062556575a2878d7e197400000000000000000000000000000000000000000000000000000000000000000000000000000000021e21a3668134f6072ba6624aa7064bd5076a8ea000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004a73219fbcbeb2f0bc4c01690800000000000000000006ae718916430000a0062556575a2878d7e197400000000000000000000000000000000000000000000000000000000000000000000000000000000021e21a3668134f6072ba6624aa7064bd5076a8ea00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
parameter UDP_BIT_PHV_SEG_02  = 4096'h5860481e6a3e240908b57e840800000000000000000005bc2637025b00006c11078364a10cced39c4e31000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d981000069aa4a5400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005860481e6a3e240908b57e840800000000000000000005bc2637025b00006c11078364a10cced39c4e31000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d981000069aa4a540000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


reg result_correct_SEG_02 = 1'b0 ;
reg [4095:0] data_temp_icmp_SEG_02 = 'b0 ;
reg [4095:0] data_temp_tcp_SEG_02  = 'b0 ;
reg [4095:0] data_temp_udp_SEG_02  = 'b0 ;
wire [4095:0] wire_data_temp_icmp_SEG_02  ;
wire [4095:0] wire_data_temp_tcp_SEG_02   ;
wire [4095:0] wire_data_temp_udp_SEG_02   ;


assign wire_data_temp_icmp_SEG_02 =  data_o&ICMP_BIT_MASK_SEG_02;
assign wire_data_temp_tcp_SEG_02  =  data_o&TCP_BIT_MASK_SEG_02;
assign wire_data_temp_udp_SEG_02  =  data_o&UDP_BIT_MASK_SEG_02;

reg flag_icmp_SEG_02 ;
reg flag_tcp_SEG_02  ;
reg flag_udp_SEG_02  ;

always @(negedge clk) begin
    // if ( dval_o == 1'b1 ) begin
        data_temp_icmp_SEG_02 <= (data_o&ICMP_BIT_MASK_SEG_02)^ICMP_BIT_PHV_SEG_02    ;
        data_temp_tcp_SEG_02  <= (data_o&TCP_BIT_MASK_SEG_02 )^TCP_BIT_PHV_SEG_02     ;
        data_temp_udp_SEG_02  <= (data_o&UDP_BIT_MASK_SEG_02 )^UDP_BIT_PHV_SEG_02     ;
        
        flag_icmp_SEG_02 <=  ((data_o&ICMP_BIT_MASK_SEG_02) == ICMP_BIT_PHV_SEG_02); // |((data_o&ICMP_BIT_MASK)^ICMP_BIT_PHV ) ;
        flag_tcp_SEG_02  <= |((data_o&TCP_BIT_MASK_SEG_02 )^TCP_BIT_PHV_SEG_02  ) ;
        flag_udp_SEG_02  <= |((data_o&UDP_BIT_MASK_SEG_02 )^UDP_BIT_PHV_SEG_02  ) ;


        if ( !((data_o&ICMP_BIT_MASK_SEG_02)^ICMP_BIT_PHV_SEG_02) ) begin // data_o&ICMP_BIT_MASK == ICMP_BIT_PHV
            result_correct_SEG_02 <= 1'b1;
        end
        else if (!((data_o&TCP_BIT_MASK_SEG_02 )^TCP_BIT_PHV_SEG_02)) begin // data_o&TCP_BIT_MASK == TCP_BIT_PHV
            result_correct_SEG_02 <= 1'b1;
        end
        else if(!((data_o&UDP_BIT_MASK_SEG_02 )^UDP_BIT_PHV_SEG_02)) begin // data_o&UDP_BIT_MASK == UDP_BIT_PHV
            result_correct_SEG_02 <= 1'b1;
        end
        else begin
            result_correct_SEG_02 <= 1'b0;
        end
    // end
end



parameter ICMP_BIT_MASK_SEG_04 = 4096'hffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffff0000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffff0000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffff0000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffff0000000000000000000000000000;
parameter TCP_BIT_MASK_SEG_04  = 4096'hffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000;
parameter UDP_BIT_MASK_SEG_04  = 4096'hffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffff000000000000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffff000000000000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffff000000000000000000000000000000000000ffffffffffffffffffffffffffff0000000000000000ffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffff000000000000000000000000000000000000;


parameter ICMP_BIT_PHV_SEG_04 = 4096'heed6640c13fe75b83ed539a908000000000000000000057ce2d64b9b0000d80105f530670ec2cc885628000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008d026080000000000000000000000000000eed6640c13fe75b83ed539a908000000000000000000057ce2d64b9b0000d80105f530670ec2cc885628000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008d026080000000000000000000000000000eed6640c13fe75b83ed539a908000000000000000000057ce2d64b9b0000d80105f530670ec2cc885628000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008d026080000000000000000000000000000eed6640c13fe75b83ed539a908000000000000000000057ce2d64b9b0000d80105f530670ec2cc885628000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008d026080000000000000000000000000000;
parameter TCP_BIT_PHV_SEG_04  = 4096'h4a73219fbcbeb2f0bc4c01690800000000000000000006ae718916430000a0062556575a2878d7e197400000000000000000000000000000000000000000000000000000000000000000000000000000000021e21a3668134f6072ba6624aa7064bd5076a8ea00000000000000000000000000000000000000000000000000004a73219fbcbeb2f0bc4c01690800000000000000000006ae718916430000a0062556575a2878d7e197400000000000000000000000000000000000000000000000000000000000000000000000000000000021e21a3668134f6072ba6624aa7064bd5076a8ea00000000000000000000000000000000000000000000000000004a73219fbcbeb2f0bc4c01690800000000000000000006ae718916430000a0062556575a2878d7e197400000000000000000000000000000000000000000000000000000000000000000000000000000000021e21a3668134f6072ba6624aa7064bd5076a8ea00000000000000000000000000000000000000000000000000004a73219fbcbeb2f0bc4c01690800000000000000000006ae718916430000a0062556575a2878d7e197400000000000000000000000000000000000000000000000000000000000000000000000000000000021e21a3668134f6072ba6624aa7064bd5076a8ea0000000000000000000000000000000000000000000000000000;
parameter UDP_BIT_PHV_SEG_04  = 4096'h5860481e6a3e240908b57e840800000000000000000005bc2637025b00006c11078364a10cced39c4e31000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d981000069aa4a540000000000000000000000000000000000005860481e6a3e240908b57e840800000000000000000005bc2637025b00006c11078364a10cced39c4e31000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d981000069aa4a540000000000000000000000000000000000005860481e6a3e240908b57e840800000000000000000005bc2637025b00006c11078364a10cced39c4e31000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d981000069aa4a540000000000000000000000000000000000005860481e6a3e240908b57e840800000000000000000005bc2637025b00006c11078364a10cced39c4e31000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d981000069aa4a54000000000000000000000000000000000000;


reg result_correct_SEG_04 = 1'b0 ;
reg [4095:0] data_temp_icmp_SEG_04 = 'b0 ;
reg [4095:0] data_temp_tcp_SEG_04  = 'b0 ;
reg [4095:0] data_temp_udp_SEG_04  = 'b0 ;
wire [4095:0] wire_data_temp_icmp_SEG_04  ;
wire [4095:0] wire_data_temp_tcp_SEG_04   ;
wire [4095:0] wire_data_temp_udp_SEG_04   ;


assign wire_data_temp_icmp_SEG_04 =  data_o&ICMP_BIT_MASK_SEG_04;
assign wire_data_temp_tcp_SEG_04  =  data_o&TCP_BIT_MASK_SEG_04;
assign wire_data_temp_udp_SEG_04  =  data_o&UDP_BIT_MASK_SEG_04;

reg flag_icmp_SEG_04 ;
reg flag_tcp_SEG_04  ;
reg flag_udp_SEG_04  ;

always @(negedge clk) begin
    // if ( dval_o == 1'b1 ) begin
        data_temp_icmp_SEG_04 <= (data_o&ICMP_BIT_MASK_SEG_04)^ICMP_BIT_PHV_SEG_04    ;
        data_temp_tcp_SEG_04  <= (data_o&TCP_BIT_MASK_SEG_04 )^TCP_BIT_PHV_SEG_04     ;
        data_temp_udp_SEG_04  <= (data_o&UDP_BIT_MASK_SEG_04 )^UDP_BIT_PHV_SEG_04     ;
        
        flag_icmp_SEG_04 <=  ((data_o&ICMP_BIT_MASK_SEG_04) == ICMP_BIT_PHV_SEG_04); // |((data_o&ICMP_BIT_MASK)^ICMP_BIT_PHV ) ;
        flag_tcp_SEG_04  <= |((data_o&TCP_BIT_MASK_SEG_04 )^TCP_BIT_PHV_SEG_04  ) ;
        flag_udp_SEG_04  <= |((data_o&UDP_BIT_MASK_SEG_04 )^UDP_BIT_PHV_SEG_04  ) ;


        if ( !((data_o&ICMP_BIT_MASK_SEG_04)^ICMP_BIT_PHV_SEG_04) ) begin // data_o&ICMP_BIT_MASK == ICMP_BIT_PHV
            result_correct_SEG_04 <= 1'b1;
        end
        else if (!((data_o&TCP_BIT_MASK_SEG_04 )^TCP_BIT_PHV_SEG_04)) begin // data_o&TCP_BIT_MASK == TCP_BIT_PHV
            result_correct_SEG_04 <= 1'b1;
        end
        else if(!((data_o&UDP_BIT_MASK_SEG_04 )^UDP_BIT_PHV_SEG_04)) begin // data_o&UDP_BIT_MASK == UDP_BIT_PHV
            result_correct_SEG_04 <= 1'b1;
        end
        else begin
            result_correct_SEG_04 <= 1'b0;
        end
    // end
end






// always @(negedge clk) begin
//     // if ( dval_o == 1'b1 ) begin
//         data_temp_icmp <= (data_o&ICMP_BIT_MASK)^ICMP_BIT_PHV    ;
//         data_temp_tcp  <= (data_o&TCP_BIT_MASK )^TCP_BIT_PHV     ;
//         data_temp_udp  <= (data_o&UDP_BIT_MASK )^UDP_BIT_PHV     ;
        
//         flag_icmp <=  ((data_o&ICMP_BIT_MASK) == ICMP_BIT_PHV); // |((data_o&ICMP_BIT_MASK)^ICMP_BIT_PHV ) ;
//         flag_tcp  <= |((data_o&TCP_BIT_MASK )^TCP_BIT_PHV  ) ;
//         flag_udp  <= |((data_o&UDP_BIT_MASK )^UDP_BIT_PHV  ) ;


//         if ( !((data_o&ICMP_BIT_MASK)^ICMP_BIT_PHV) ) begin // data_o&ICMP_BIT_MASK == ICMP_BIT_PHV
//             result_correct <= 1'b1;
//         end
//         else if (!((data_o&TCP_BIT_MASK )^TCP_BIT_PHV)) begin // data_o&TCP_BIT_MASK == TCP_BIT_PHV
//             result_correct <= 1'b1;
//         end
//         else if(!((data_o&UDP_BIT_MASK )^UDP_BIT_PHV)) begin // data_o&UDP_BIT_MASK == UDP_BIT_PHV
//             result_correct <= 1'b1;
//         end
//         else begin
//             result_correct <= 1'b0;
//         end
//     // end
// end



endmodule


















// test_pex_ibf_pdep_bf_top #(
//     .DATA_WIDTH ( DATA_WIDTH )
    
//     )
//  u_test_pex_ibf_pdep_bf_top (
//     .clk                     ( clk                                       ),
//     .rst                     ( rst                                       ),
//     .mode_i                  ( mode_i            [MODE_WIDTH-1:0]        ),
//     .dval_i                  ( dval_i                                    ),
//     .data_i                  ( data_i            [DATA_WIDTH-1:0]        ),
//     .ibf_sram_sel_2_2        ( ibf_sram_sel_2_2  [7:0]                   ),
//     .ibf_wr_en_2_2           ( ibf_wr_en_2_2                             ),
//     .ibf_wr_cfg_2_2          ( ibf_wr_cfg_2_2    [IBF_CFG_WIDTH_2_2-1:0] ),
//     .ibf_wr_en_2_1           ( ibf_wr_en_2_1                             ),
//     .ibf_wr_cfg_2_1          ( ibf_wr_cfg_2_1    [IBF_CFG_WIDTH_2_1-1:0] ),
//     .bf_sram_sel_2_2         ( bf_sram_sel_2_2   [7:0]                   ),
//     .bf_wr_en_2_2            ( bf_wr_en_2_2                              ),
//     .bf_wr_cfg_2_2           ( bf_wr_cfg_2_2     [BF_CFG_WIDTH_2_2-1:0]  ),

//     .dval_o                  ( dval_o                                    ),
//     .data_o                  ( data_o            [DATA_WIDTH-1:0]        )
// );
